module FSM();
endmodule